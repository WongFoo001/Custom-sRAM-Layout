magic
tech sky130A
timestamp 1647623508
<< nwell >>
rect -265 50 -119 145
rect -344 -34 -119 50
rect -265 -114 -119 -34
<< nsubdiff >>
rect -316 9 -267 17
rect -316 -9 -302 9
rect -283 -9 -267 9
rect -316 -15 -267 -9
<< nsubdiffcont >>
rect -302 -9 -283 9
<< poly >>
rect -448 108 -137 124
rect -424 -35 -406 108
rect -195 -35 -177 108
rect -424 -44 -177 -35
rect -424 -50 -302 -44
rect -424 -70 -406 -50
rect -450 -85 -406 -70
rect -330 -69 -302 -50
rect -276 -50 -177 -44
rect -276 -69 -249 -50
rect -330 -77 -249 -69
rect -195 -70 -177 -50
rect -195 -85 -138 -70
<< polycont >>
rect -302 -69 -276 -44
<< locali >>
rect -321 92 -259 102
rect -321 72 -299 92
rect -280 72 -259 92
rect -321 33 -259 72
rect -348 9 -227 33
rect -348 -9 -302 9
rect -283 -9 -227 9
rect -348 -18 -227 -9
rect -330 -44 -249 -40
rect -330 -69 -302 -44
rect -276 -69 -249 -44
<< viali >>
rect -299 72 -280 92
rect -300 -68 -278 -45
<< metal1 >>
rect -448 -111 -407 148
rect -366 -78 -325 150
rect -309 111 -266 114
rect -309 110 -302 111
rect -310 83 -302 110
rect -272 83 -266 111
rect -310 72 -299 83
rect -280 72 -266 83
rect -310 67 -266 72
rect -367 -112 -325 -78
rect -305 -45 -273 -37
rect -305 -68 -300 -45
rect -278 -68 -273 -45
rect -305 -84 -273 -68
rect -244 -114 -203 151
rect -176 -114 -135 151
<< via1 >>
rect -302 92 -272 111
rect -302 83 -299 92
rect -299 83 -280 92
rect -280 83 -272 92
<< metal2 >>
rect -448 111 -137 115
rect -448 83 -302 111
rect -272 83 -137 111
rect -448 81 -137 83
rect -448 3 -138 37
rect -448 -80 -138 -46
<< labels >>
rlabel locali -290 45 -290 45 1 VPB
<< end >>
