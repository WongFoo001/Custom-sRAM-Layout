magic
tech sky130A
timestamp 1647646066
<< pwell >>
rect -335 157 -249 158
rect -337 -2 -236 139
<< psubdiff >>
rect -310 116 -270 134
rect -310 99 -299 116
rect -282 99 -270 116
rect -310 80 -270 99
rect -310 63 -299 80
rect -282 63 -270 80
rect -310 48 -270 63
<< psubdiffcont >>
rect -299 99 -282 116
rect -299 63 -282 80
<< poly >>
rect -448 151 -137 166
rect -348 -5 -330 151
rect -249 -5 -231 151
rect -348 -14 -231 -5
rect -348 -28 -300 -14
rect -448 -36 -300 -28
rect -278 -28 -231 -14
rect -278 -36 -138 -28
rect -448 -43 -138 -36
rect -448 -44 -313 -43
<< polycont >>
rect -300 -36 -278 -14
<< locali >>
rect -321 116 -259 145
rect -321 99 -299 116
rect -282 99 -259 116
rect -321 80 -259 99
rect -321 79 -299 80
rect -282 79 -259 80
rect -321 56 -300 79
rect -278 56 -259 79
rect -321 41 -259 56
rect -330 -36 -300 -5
rect -278 -36 -249 -5
rect -330 -43 -249 -36
<< viali >>
rect -300 63 -299 79
rect -299 63 -282 79
rect -282 63 -278 79
rect -300 56 -278 63
rect -300 -14 -278 -2
rect -300 -25 -278 -14
<< metal1 >>
rect -448 -72 -407 194
rect -381 -72 -340 194
rect -308 79 -270 96
rect -308 51 -302 79
rect -276 51 -270 79
rect -308 46 -270 51
rect -305 -2 -273 6
rect -305 -25 -300 -2
rect -278 -25 -273 -2
rect -305 -41 -273 -25
rect -244 -72 -203 194
rect -176 -72 -135 194
<< via1 >>
rect -302 56 -300 79
rect -300 56 -278 79
rect -278 56 -276 79
rect -302 51 -276 56
<< metal2 >>
rect -448 124 -137 158
rect -448 79 -138 80
rect -448 51 -302 79
rect -276 51 -138 79
rect -448 46 -138 51
rect -448 -37 -138 -3
<< labels >>
rlabel locali -289 90 -289 90 1 VNB
<< end >>
