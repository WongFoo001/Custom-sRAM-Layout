magic
tech sky130A
magscale 1 2
timestamp 1647621430
<< nwell >>
rect 118 -142 410 388
<< nmos >>
rect -122 302 -38 332
rect -122 156 -38 186
rect -122 60 -38 90
rect -122 -86 -38 -56
<< pmos >>
rect 170 156 254 186
rect 170 60 254 90
<< ndiff >>
rect -122 378 -38 388
rect -122 344 -98 378
rect -64 344 -38 378
rect -122 332 -38 344
rect -122 280 -38 302
rect -122 246 -96 280
rect -62 246 -38 280
rect -122 186 -38 246
rect -238 140 -176 154
rect -238 106 -225 140
rect -191 138 -176 140
rect -122 138 -38 156
rect -191 106 -38 138
rect -238 94 -176 106
rect -122 90 -38 106
rect -122 0 -38 60
rect -122 -34 -98 0
rect -64 -34 -38 0
rect -122 -56 -38 -34
rect -122 -98 -38 -86
rect -122 -132 -98 -98
rect -64 -132 -38 -98
rect -122 -142 -38 -132
<< pdiff >>
rect 170 278 254 286
rect 170 244 196 278
rect 230 244 254 278
rect 170 186 254 244
rect 170 140 254 156
rect 308 142 372 152
rect 308 140 326 142
rect 170 108 326 140
rect 360 108 372 142
rect 170 90 254 108
rect 308 98 372 108
rect 170 2 254 60
rect 170 -8 196 2
rect 168 -32 196 -8
rect 230 -32 254 2
rect 168 -40 254 -32
<< ndiffc >>
rect -98 344 -64 378
rect -96 246 -62 280
rect -225 106 -191 140
rect -98 -34 -64 0
rect -98 -132 -64 -98
<< pdiffc >>
rect 196 244 230 278
rect 326 108 360 142
rect 196 -32 230 2
<< poly >>
rect -246 302 -122 332
rect -38 302 378 332
rect -2 200 122 210
rect -2 186 24 200
rect -150 156 -122 186
rect -38 166 24 186
rect 66 186 122 200
rect 66 166 170 186
rect -38 156 170 166
rect 254 156 292 186
rect -150 60 -122 90
rect -38 80 170 90
rect -38 60 60 80
rect 0 46 60 60
rect 102 60 170 80
rect 254 60 292 90
rect 102 46 122 60
rect 0 34 122 46
rect -248 -86 -122 -56
rect -38 -86 378 -56
<< polycont >>
rect 24 166 66 200
rect 60 46 102 80
<< locali >>
rect -150 384 290 388
rect -150 378 -52 384
rect -150 344 -98 378
rect -64 350 -52 378
rect -18 350 290 384
rect -64 344 290 350
rect -150 342 290 344
rect -122 280 254 284
rect -122 246 -96 280
rect -62 278 254 280
rect -62 246 196 278
rect -122 244 196 246
rect 230 244 254 278
rect -122 242 254 244
rect -38 200 86 208
rect -38 166 24 200
rect 66 166 86 200
rect -248 140 -170 160
rect -248 106 -225 140
rect -191 106 -170 140
rect -248 90 -170 106
rect -38 156 86 166
rect -38 4 -2 156
rect 120 90 160 242
rect 302 142 380 160
rect 302 108 326 142
rect 360 108 380 142
rect 302 90 380 108
rect 38 80 160 90
rect 38 46 60 80
rect 102 46 160 80
rect 38 38 160 46
rect -122 2 254 4
rect -122 0 196 2
rect -122 -34 -98 0
rect -64 -32 196 0
rect 230 -32 254 2
rect -64 -34 254 -32
rect -122 -38 254 -34
rect -150 -98 290 -96
rect -150 -132 -98 -98
rect -64 -102 290 -98
rect -64 -132 184 -102
rect -150 -136 184 -132
rect 220 -136 290 -102
rect -150 -142 290 -136
<< viali >>
rect -52 350 -18 384
rect -225 106 -191 140
rect 326 108 360 142
rect 184 -136 220 -102
<< metal1 >>
rect -248 150 -166 388
rect -248 96 -236 150
rect -180 96 -166 150
rect -248 -144 -166 96
rect -84 384 -2 390
rect -84 350 -52 384
rect -18 350 -2 384
rect -84 -144 -2 350
rect 160 -102 242 390
rect 160 -136 184 -102
rect 220 -136 242 -102
rect 160 -142 242 -136
rect 296 306 378 388
rect 296 252 317 306
rect 369 252 378 306
rect 296 142 378 252
rect 296 108 326 142
rect 360 108 378 142
rect 160 -144 240 -142
rect 296 -144 378 108
<< via1 >>
rect -236 140 -180 150
rect -236 106 -225 140
rect -225 106 -191 140
rect -191 106 -180 140
rect -236 96 -180 106
rect 317 252 369 306
<< metal2 >>
rect -244 314 -120 316
rect -244 306 378 314
rect -244 252 317 306
rect 369 252 378 306
rect -244 248 378 252
rect -246 150 378 158
rect -246 96 -236 150
rect -180 96 378 150
rect -246 92 378 96
rect -246 -72 372 -6
<< labels >>
rlabel locali -6 366 -6 366 1 BL
port 4 n
rlabel locali 148 -122 148 -122 1 BR
port 5 n
rlabel metal1 338 196 338 196 1 vdd
rlabel poly 60 324 60 324 1 WL
rlabel poly 70 -78 70 -78 1 WL
rlabel locali 56 246 56 246 1 Q
rlabel locali 70 0 70 0 1 QB
rlabel metal2 -204 -38 -204 -38 1 WL
rlabel metal1 -200 202 -200 202 1 gnd
<< end >>
