* NGSPICE file created from cell_1rw.ext - technology: sky130A

.subckt cell_1rw BL BR VSUBS w_130_n80#
X0 BL WL Q VSUBS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=2.436e+11p ps=2e+06u w=420000u l=150000u
X1 gnd Q QB VSUBS sky130_fd_pr__nfet_01v8 ad=2.655e+11p pd=2.88e+06u as=2.436e+11p ps=2e+06u w=420000u l=150000u
X2 QB WL BR VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X3 Q QB gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 vdd Q QB w_130_n80# sky130_fd_pr__pfet_01v8 ad=2.682e+11p pd=2.9e+06u as=2.116e+11p ps=1.86e+06u w=420000u l=150000u
X5 Q QB vdd w_130_n80# sky130_fd_pr__pfet_01v8 ad=2.1e+11p pd=1.84e+06u as=0p ps=0u w=420000u l=150000u
.ends

